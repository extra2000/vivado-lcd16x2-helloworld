`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////////////////////
//234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567
//        1         2         3         4         5         6         7         8         9
//------------------------------------------------------------------------------------------------
// 8MHz clock generator test bench
//////////////////////////////////////////////////////////////////////////////////////////////////


module clock_generator_8mhz_tb;

  reg  clk_i = 0;
  wire clk_o;

  clock_generator_8mhz UUT(
    .clk_i(clk_i),
    .clk_o(clk_o)
  );

  // Delaying 8ns before inverting r_clock to simulate 125MHz clock.
  always #8 clk_i <= !clk_i;

endmodule
